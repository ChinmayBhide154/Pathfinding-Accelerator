module Pathfinding (
    input logic temp1,
    output logic temp2
);
    
    
endmodule