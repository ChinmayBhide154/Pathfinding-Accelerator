//===================================================================
// Design name:		Parameters for Floating Point Unit DD192
// Note: 			Addition, Subtraction, Multiply, Divide, Square Root
// Project name:	A 32 bit single precision Floating Point Unit DD192 
// Author:			hungbk99
//===================================================================

package	FPU_192_Package;
	
	parameter	FORMAT_LENGTH = 32;
	parameter	EXPONENT_LENGTH = 8;
	parameter	FRACTION_LENGTH = 23;
	parameter 	NORMALIZE_MANTISSA_LENGTH = 24;
	parameter 	DIVIDEND_LENGTH = 24;
	parameter 	DIVISOR_LENGTH = 24;
	parameter	QUOTIENT_LENGTH = 24;

endpackage
