module CoordinateCollector (
    input logic reset,
    input logic clk,
    input logic [255:0] xCoord,
    input logic [255:0] yCoord,
    input logic transition,
    input logic enterNewCoord,
    input logic finishInit,

    output logic done
);


typedef enum logic [1:0] {  
    GET_X = 2'b00,
    GET_Y = 2'b01,
    UPDATE_MEM = 2'b10,
    FINISH = 2'b11
} stateType;

stateType state = GET_X;

logic [1:0] next;

always_ff @(posedge clk or posedge reset) begin
    if(reset) state <= GET_X;
    else state <= next;
end

always_comb begin
    case(state)
        GET_X: if(transition) next = GET_Y;
                else next = GET_X;

        GET_Y: if(transition) next = UPDATE_MEM;
                else next = GET_Y;

        UPDATE_MEM: if(enterNewCoord) next = GET_X;
                    else if(finishInit) next = FINISH;
                    else next = UPDATE_MEM;

        FINISH: next = FINISH;
    endcase
end


endmodule
